* SPICE netlist written by S-Edit Win32 6.00
* Written on Mar 28, 2024 at 19:34:30

* Waveform probing commands
.probe
.options probefilename="DFF"
+ probesdbfile="C:\Users\IDEAL\Desktop\CA1\part 2\DFF.sdb"
+ probetopmodule="ShR4bit"

* No Ports in cell: PageID_Tanner
* End of module with no ports: PageID_Tanner

.SUBCKT Pad_Bond SIGNAL Subs
C1 SIGNAL Subs 0.25pF
* Page Size:  5x7
* S-Edit  Output Pad
* Designed by: D.Gunawan, J.Luo, K.Schaefer  Mar 28, 2024  11:21:00
* Schematic generated by S-Edit
* from file C:\Users\IDEAL\Desktop\CA1\part 2\DFF / module Pad_Bond / page Page0 
.ENDS

.SUBCKT PadBidirHE_2.0u DataIn DataInB DataInUnBuf DataOut OE Pad Gnd Subs Vdd
MN_4_1 OEB OE Gnd Gnd NMOS W=22u L=2u AS=66p AD=66p PS=24u PD=24u M=1
MN_4_2 N29 DataOut Gnd Gnd NMOS W=22u L=2u AS=66p AD=66p PS=24u PD=24u M=1
MN_4_3 N20 OE N29 Gnd NMOS W=22u L=2u AS=66p AD=66p PS=24u PD=24u M=1
MN_4_4 N29 OEB Gnd Gnd NMOS W=22u L=2u AS=66p AD=66p PS=24u PD=24u M=1
MN_4_5 Pad N29 Gnd Gnd NMOS W=22u L=2u AS=66p AD=66p PS=24u PD=24u M=10
MN_4_6 DataInB DataInUnBuf Gnd Gnd NMOS W=22u L=2u AS=66p AD=66p PS=24u PD=24u M=2
MN_4_7 DataIn DataInB Gnd Gnd NMOS W=22u L=2u AS=66p AD=66p PS=24u PD=24u M=4
XPad_Bond_1 Pad Subs Pad_Bond
* Page Size:  5x7
* S-Edit  Bidirectional Pad
* Designed by: D.Gunawan, J.Luo  Mar 28, 2024  11:21:00
* Schematic generated by S-Edit
* from file C:\Users\IDEAL\Desktop\CA1\part 2\DFF / module PadBidirHE_2.0u / page Page0 
MP_4_1 OEB OE Vdd Vdd PMOS W=22u L=2u AS=66p AD=66p PS=24u PD=24u M=1
MP_4_2 N20 DataOut Vdd Vdd PMOS W=22u L=2u AS=66p AD=66p PS=24u PD=24u M=2
MP_4_3 N29 OEB N20 Vdd PMOS W=22u L=2u AS=66p AD=66p PS=24u PD=24u M=2
MP_4_4 N20 OE Vdd Vdd PMOS W=22u L=2u AS=66p AD=66p PS=24u PD=24u M=1
MP_4_5 Pad N20 Vdd Vdd PMOS W=22u L=2u AS=66p AD=66p PS=24u PD=24u M=10
MP_4_6 DataInB DataInUnBuf Vdd Vdd PMOS W=22u L=2u AS=66p AD=66p PS=24u PD=24u M=2
MP_4_7 DataIn DataInB Vdd Vdd PMOS W=22u L=2u AS=66p AD=66p PS=24u PD=24u M=4
R1 Pad DataInUnBuf 100 TC1=0.0 TC2=0.0
.ENDS

.SUBCKT PadBidirHE DataIn DataInB DataInUnBuf DataOut OE Pad Gnd Subs Vdd
XPadBidirHE_2.0u_1 DataIn DataInB DataInUnBuf DataOut OE Pad Gnd Subs Vdd
+ PadBidirHE_2.0u
* Page Size:  5x7
* S-Edit  Bidirectional Pad
* Designed by: D.Gunawan, J.Luo  Mar 28, 2024  11:21:00
* Schematic generated by S-Edit
* from file C:\Users\IDEAL\Desktop\CA1\part 2\DFF / module PadBidirHE / page Page0 
.ENDS

.SUBCKT PadOut DataOut Pad Gnd Subs Vdd
XPadBidirHE_1 N6 N5 N4 DataOut Vdd Pad Gnd Subs Vdd PadBidirHE
* Page Size:  5x7
* S-Edit  Output Pad
* Designed by: D.Gunawan, J.Luo  Mar 28, 2024  11:21:00
* Schematic generated by S-Edit
* from file C:\Users\IDEAL\Desktop\CA1\part 2\DFF / module PadOut / page Page0 
.ENDS

.SUBCKT PadInC DataIn DataInB DataInUnBuf Pad Gnd Subs Vdd
XPadBidirHE_1 DataIn DataInB DataInUnBuf Gnd Gnd Pad Gnd Subs Vdd PadBidirHE
* Page Size:  5x7
* S-Edit  Input Pad
* Designed by: D.Gunawan, J.Luo  Mar 28, 2024  11:19:10
* Schematic generated by S-Edit
* from file C:\Users\IDEAL\Desktop\CA1\part 2\DFF / module PadInC / page Page0 
.ENDS

.SUBCKT NAND2 A B Out Gnd Vdd
M3 Out B 1 Gnd NMOS W='28*l' L='2*l' AS='148*l*l' AD='84*l*l' PS='68*l' PD='34*l' M=1
M4 1 A Gnd Gnd NMOS W='28*l' L='2*l' AS='84*l*l' AD='144*l*l' PS='34*l' PD='68*l' M=1
* Page Size:  5x7
* S-Edit  2-Input NAND Gate (TIB)
* Designed by: J. Luo  Mar 28, 2024  11:17:13
* Schematic generated by S-Edit
* from file C:\Users\IDEAL\Desktop\CA1\part 2\DFF / module NAND2 / page Page0 
M2 Out B Vdd Vdd PMOS W='28*l' L='2*l' AS='144*l*l' AD='84*l*l' PS='68*l' PD='34*l' M=1
M1 Out A Vdd Vdd PMOS W='28*l' L='2*l' AS='84*l*l' AD='144*l*l' PS='34*l' PD='68*l' M=1
.ENDS

.SUBCKT Inv A Out Gnd Vdd
M2 Out A Gnd Gnd NMOS W='28*l' L='2*l' AS='148*l*l' AD='144*l*l' PS='68*l' PD='68*l' M=1
* Page Size:  5x7
* S-Edit  Inverter (TIB)
* Designed by: J. Luo  Mar 28, 2024  11:17:13
* Schematic generated by S-Edit
* from file C:\Users\IDEAL\Desktop\CA1\part 2\DFF / module Inv / page Page0 
M1 Out A Vdd Vdd PMOS W='28*l' L='2*l' AS='148*l*l' AD='144*l*l' PS='68*l' PD='68*l' M=1
.ENDS

.SUBCKT DFF Clk D Q Qbar Gnd Vdd
XInv_1 Clk N8 Gnd Vdd Inv
XInv_2 D N2 Gnd Vdd Inv
XNAND2_1 D Clk N5 Gnd Vdd NAND2
XNAND2_2 Clk N2 N4 Gnd Vdd NAND2
XNAND2_3 N6 N4 N7 Gnd Vdd NAND2
XNAND2_4 N5 N7 N6 Gnd Vdd NAND2
XNAND2_5 N6 N8 N10 Gnd Vdd NAND2
XNAND2_6 N8 N7 N9 Gnd Vdd NAND2
XNAND2_7 Q N9 Qbar Gnd Vdd NAND2
XNAND2_8 N10 Qbar Q Gnd Vdd NAND2
.ENDS

* Main circuit: ShR4bit
XDFF_1 N2 N1 N5 N4 Gnd Vdd DFF
XDFF_3 N2 N5 N9 N8 Gnd Vdd DFF
XDFF_4 N2 N9 N13 N12 Gnd Vdd DFF
XDFF_5 N2 N13 N15 N16 Gnd Vdd DFF
XPadInC_1 N1 N11 N7 Serial_Input Gnd Subs Vdd PadInC
XPadInC_2 N2 N19 N18 Clk Gnd Subs Vdd PadInC
XPadOut_1 N15 Serial_Output Gnd Subs Vdd PadOut
* End of main circuit: ShR4bit

***********library*************
.inc 0.5micron.lib
*******************************
.PARAM l = 0.5u

*************Inputs************
Vpulse Clk 0 PULSE(0 5 0 1ps 1ps 50ns 100ns)
VserIn Serial_Input 0 DC 0
*******************************



*******************************
.op
.tran 1ns 2us
.options post=2
.measure tran power_avg AVG power from=0n to=160n
*******************************

